package my_package;
  parameter ROWS = 4;
  parameter COLUMNS = 4;
  parameter PAKG_SIZE = 32;
  parameter FIFO_DEPTH = 10;
endpackage
