`define PAKG_SIZE 38
`define FIFO_DEPTH 3
